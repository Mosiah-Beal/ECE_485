package my_struct_package;


// define MESI states
typedef enum logic [1:0] {
	I = 2'b00, // Invalid
	S = 2'b01, // Shared
	E = 2'b10, // Exclusive
	M = 2'b11  // Modified
} states_t;

// Address struct, unpacks 32-bit address into tag, set index, and byte offset
typedef struct packed {
	logic [11:0] tag;         // 12 bits for tag
	logic [13:0] set_index;   // 14 bits for set index
	logic [5:0]  byte_offset; // 6 bits for byte offset
} address_t;

// Processor instruction struct, contains instruction, address, and processor ID
typedef struct packed {
    logic [3:0] n;             // instruction
    address_t address;      // 32-bit address
} command_t;

// Cache line struct, contains tag, LRU, MESI bits, and data
typedef struct packed {
	logic [11:0] tag;         // 12 bits for tag
	logic [2:0] LRU;          // 3 bits for LRU
	states_t MESI_bits;    // 2 bits for MESI states
	logic [31:0] data;        // 512 bits for data
} cache_line_t;



endpackage

