module mesi_ctrl();

endmodule
